** sch_path: /home/cmaier/EDA/efabless/chipalooza2024/sky130_rodovalho_ip__lpopamp/cace/tb_lpopamp_open_op.sch
**.subckt tb_lpopamp_open_op
Xdut out ip out avdd avss en enb ibias sky130_rodovalho_ip__lpopamp
v_avss GND net1 0
v_avdd avdd net1 dc 3.3
v_en en avss 3.3
v_enb enb avss 0
i_ibias avdd ibias xibias
c_l out avss {xcl} m=1
v_ip ip avss dc xvin
**** begin user architecture code


.param mc_mm_switch=0
.temp 25




.option gmin=1e-12
.option rshunt=1e12
.control
  op
  let idd = op.i(v_avdd)
  set wr_singlescale
  wrdata ngspice/idd_1.data idd
  quit
.endc




.param xavdd  = 3.3
.param xvin   = 1.65

.param xibias = 10u
.param xcl    = 30p



** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130A/libs.tech/combined/sky130.lib.spice tt


**** end user architecture code
**.ends
.GLOBAL GND
.end
